-------------------------------------------------------------------------------
-- Title      : Trigger Hold
-- Project    : Source files in two directories, custom library name, VHDL'87
-------------------------------------------------------------------------------
-- File       : st_comb.vhd
-- Author     :   <kimei@fyspc-epf02>
-- Company    : 
-- Created    : 2011-03-15
-- Last update: 2011-03-17
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: Synchronous trigger part of the CTU in COMPET
-------------------------------------------------------------------------------
-- Copyright (c) 2011 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2011-03-08  1.0      kimei   Created
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

library work;
use work.components.all;
use work.constants.all;
use work.functions.all;

entity trigger_hold is
  port (
    edge_in_b : in  std_logic;
    mclk      : in  std_logic;
    rst_b     : in  std_logic;
    trig_hold : out std_logic);
end trigger_hold;


architecture comb of trigger_hold is
  signal counter : integer range 15 downto 0;
  
begin 
  hold_signal: process (mclk, rst_b, edge_in_b)
  begin  -- process hold_signal
    if rst_b = '0' then                 
      trig_hold <= '0';
      counter <= 0;
    elsif edge_in_b = '0' and counter = 0 then
      counter <= 1;
    elsif mclk'event and mclk = '1' then
      if counter /= 0 then
        trig_hold <= '1';
        counter <=  counter + 1;
      end if;

      if counter = 4 then
        counter <=  0;
        trig_hold <= '0';
      end if;
      
    end if;
  end process hold_signal;

end comb;
