-------------------------------------------------------------------------------
-- Title      : Sync Trigger
-- Project    : Source files in two directories, custom library name, VHDL'87
-------------------------------------------------------------------------------
-- File       : Sync_trigger.vhd
-- Author     :   <kimei@fyspc-epf02>
-- Company    : 
-- Created    : 2011-03-08
-- Last update: 2011-03-18
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: Synchronous trigger part of the CTU in COMPET
-------------------------------------------------------------------------------
-- Copyright (c) 2011 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2011-03-08  1.0      kimei   Created
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use ieee.numeric_std.all;     --! Numeric/arithmetical logic (IEEE standard)

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

library work;
use work.components.all;
use work.constants.all;
use work.functions.all;

entity sync_trigger is
  port (
    rst_b         : in  std_logic;
    mclk          : in  std_logic;
    trigger_in    : in  std_logic_vector(NUMBER_OF_ROCS-1 downto 0);
    trigger_in_b  : in  std_logic_vector(NUMBER_OF_ROCS-1 downto 0);
    trigger_out   : out std_logic_vector(NUMBER_OF_MODULES-1 downto 0);
    trigger_out_b : out std_logic_vector(NUMBER_OF_MODULES-1 downto 0)
    );

end sync_trigger;


architecture Behavioral of sync_trigger is
  
  subtype temp is std_logic_vector(1 downto 0);
  type    coincidence_arr is array(0 to NUMBER_OF_MODULES-1) of temp;

  signal hold_count : std_logic;        -- count from 0 to 1.. :)

  signal coincidence_array : coincidence_arr;
  signal coincidence_or    : std_logic_vector(NUMBER_OF_MODULES-1 downto 0);
  signal coincidence       : std_logic;
  signal coincidence_hold  : std_logic;

  signal trig_in_as : std_logic_vector(NUMBER_OF_ROCS - 1 downto 0);

  signal trig_out : std_logic_vector(NUMBER_OF_MODULES - 1 downto 0);

  signal leading_edge_module : std_logic_vector(NUMBER_OF_MODULES-1 downto 0);

  signal edge_det : std_logic_vector(NUMBER_OF_ROCS-1 downto 0);
  component edge_detect
    port (
      rst_b : in  std_logic;
      mclk  : in  std_logic;
      inp   : in  std_logic;
      outp  : out std_logic);
  end component;
  
  
begin
  trig_out <= (others => '1') when coincidence = '1' or coincidence_hold = '1' else (others => '0');
  -- coincidence_array(0) <= "10";
  -- coincidence_array(1)(0) <= '0';
  --coincidence_array <=  (others => "00");
  -- Not the slickest solution, but i doubt there will be more than four
  -- modules, and therefore this solution is sufficient..
  N : for n in 0 to NUMBER_OF_MODULES-1 generate
    N1 : if n = 0 generate
      leading_edge_module(n) <= '0' when all_zeros(edge_det(ROCS_IN_M1-1 downto 0)) = '1' else '1';
    end generate N1;

    N2 : if n = 1 generate
      leading_edge_module(n) <= '0' when all_zeros(edge_det(ROCS_IN_M1+ROCS_IN_M2-1 downto ROCS_IN_M1)) = '1' else '1';
    end generate N2;

    N3 : if n = 2 generate
      leading_edge_module(n) <= '0' when all_zeros(edge_det(ROCS_IN_M1+ROCS_IN_M2+ROCS_IN_M3-1 downto ROCS_IN_M1+ROCS_IN_M2)) = '1' else '1';
    end generate N3;

    N4 : if n = 3 generate
      leading_edge_module(n) <= '0' when all_zeros(edge_det(ROCS_IN_M1+ROCS_IN_M2+ROCS_IN_M3+ROCS_IN_M4-1 downto ROCS_IN_M1+ROCS_IN_M2+ROCS_IN_M3)) = '1' else '1';
    end generate N4;
  end generate N;

  G1 : for I in 0 to (NUMBER_OF_ROCS-1) generate
    diff_in : work.components.IBUFDS port map (
      -- diff_in : IBUFDS port map (
      I  => trigger_in(I),
      IB => trigger_in_b(I),
      O  => trig_in_as(I));
  end generate G1;

  G4 : for n in 0 to NUMBER_OF_MODULES-1 generate
    coincidence_or(n) <= coincidence_array(n)(1) or coincidence_array(n)(0);
  end generate G4;

  coincidence <= '1' when count_ones(coincidence_or) > 1 else '0';

  G2 : for I in 0 to (NUMBER_OF_MODULES-1) generate
    diff_out : work.components.OBUFDS port map (
      -- diff_out : OBUFDS port map (
      O  => trigger_out(I),
      OB => trigger_out_b(I),
      I  => trig_out(I));
  end generate G2;

  G3 : for I in 0 to NUMBER_OF_ROCS -1 generate
    edge_detect_1 : edge_detect
      port map (
        rst_b => rst_b,
        mclk  => mclk,
        inp   => trig_in_as(I),
        outp  => edge_det(I));
    -- purpose:
    load_sr_leading_edge : process (mclk, rst_b)
    begin  -- process load_sr_leading_edge
      if rst_b = '0' then
        coincidence_hold  <= '0';
        coincidence_array <= (others => "00");
        hold_count        <= '0';
      elsif mclk'event and mclk = '1' then
        L1 : for I in 0 to NUMBER_OF_MODULES -1 loop
          coincidence_array(I)(0) <= leading_edge_module(I);
          coincidence_array(I)(1) <= coincidence_array(I)(0);
        end loop L1;

      if coincidence = '1' then
          hold_count <= '1';
          coincidence_hold <= '1';
      elsif hold_count = '1' then
         hold_count <= '0';
         coincidence_hold <= '1';
      else
          coincidence_hold <= '0';

        end if;
        
      end if;
    end process load_sr_leading_edge;

  end generate;


  
end Behavioral;
