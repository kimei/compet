-------------------------------------------------------------------------------
-- Title      : Sync Trigger
-- Project    : Source files in two directories, custom library name, VHDL'87
-------------------------------------------------------------------------------
-- File       : st_fsm.vhd
-- Author     :   <kimei@fyspc-epf02>
-- Company    : 
-- Created    : 2011-03-15
-- Last update: 2011-03-17
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: Synchronous trigger part of the CTU in COMPET
-------------------------------------------------------------------------------
-- Copyright (c) 2011 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2011-03-08  1.0      kimei   Created
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

library work;
use work.components.all;
use work.constants.all;
use work.functions.all;

entity st_fsm is
  generic (
    NO_OF_MODULES : positive := 4);
  port (
    leading_edge_b : in  std_logic_vector(NO_OF_MODULES-1 downto 0);
    mclk           : in  std_logic;
    rst_b         : in  std_logic;
    trigger_out    : out std_logic_vector(NO_OF_MODULES-1 downto 0));
end st_fsm;


architecture FSM of st_fsm is
  type states is (INIT, FIRST_EDGE, SEC_EDGE, TRIG_DELAY, TRIG_OUT, UNDEF6, UNDEF7, UNDEF8);
  signal counter : integer range 15 downto 0;
  signal state : states;
  signal previous : std_logic_vector(leading_edge_b'length-1 downto 0);
  
begin  -- FSM
  
  fsm_proc: process (mclk, rst_b)
  begin  -- process fsm
    if rst_b = '0' then                -- asynchronous reset (active low)
      trigger_out <= (others => '0');
      previous <= (others => '1');
      state <=  INIT;
      counter <= 0;
    elsif mclk'event and mclk = '1' then  -- rising clock edge
      
      trigger_out <= (others => '0');
      
      case state is

        --init state is just there to remove annoying startup glitch in sim.
        when INIT =>
          state <= INIT;
          counter <= counter + 1;
          if counter = 10 then
            state <= FIRST_EDGE;
          end if;
        when FIRST_EDGE =>
          counter <= 0;
          previous <= (others => '1');
          if all_ones(leading_edge_b) = '1' then
            state <= FIRST_EDGE;
          else
            previous <= leading_edge_b;
            state <= SEC_EDGE;
          end if;
        when SEC_EDGE =>
            if leading_edge_b = previous then
              counter <= counter + 1;
              state <= SEC_EDGE;
            elsif counter = TRIGGER_HOLD-1 then
              state <=  FIRST_EDGE;
            else
              --counter <= 0;
              state <= TRIG_DELAY;
            end if;
            
        when TRIG_DELAY =>
            counter <= counter + 1;
            if counter = TRIGGER_DELAY-1 then
              trigger_out <= (others => '1');
              state <=  TRIG_OUT;
              counter <= 0;
            else
              state <=  TRIG_DELAY;
            end if;
       when TRIG_OUT =>
            if counter = TRIGGER_WINDOW_LENGTH-1 then
              counter <= 0;
              state <= FIRST_EDGE;
            else
            trigger_out <= (others => '1');
            counter <= counter + 1;
            end if;
            
             
        when others => null;
      end case;
    end if;
  end process fsm_proc;  

end FSM;
