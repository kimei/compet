--! \file
--! \brief Constant declarations.

--! Standard library
library ieee;
use ieee.std_logic_1164.all;  --! Standard logic
use ieee.numeric_std.all;     --! Numeric/arithmetical logic (IEEE standard)


--! \brief Constants
package constants is

end package constants;
